package tlul_pkg;

    

    
endpackage