package top_pkg;


    
endpackage